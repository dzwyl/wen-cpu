`timescale 1ns/1ps

module  data_mem(
    input   clk,
    input   result,
);

endmodule