module  data_mem(
    input   clk,
    input   result,
);

endmodule